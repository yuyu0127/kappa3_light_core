// @file controller.v
// @breif controller(コントローラ)
// @author Yusuke Matsunaga (松永 裕介)
//
// Copyright (C) 2019 Yusuke Matsunaga
// All rights reserved.
//
// [概要]
// データパスを制御する信号を生成する．
// フェイズは phasegen が生成するので
// このモジュールは完全な組み合わせ回路となる．
//
// [入力]
// cstate:     動作フェイズを表す4ビットの信号
// ir:         IRレジスタの値
// addr:       メモリアドレス(mem_wrbitsの生成に用いる)
// alu_out:    ALUの出力(分岐命令の条件判断に用いる)
//
// [出力]
// pc_sel:     PCの入力選択
// pc_ld:      PCの書き込み制御
// mem_sel:    メモリアドレスの入力選択
// mem_read:   メモリの読み込み制御
// mem_write:  メモリの書き込み制御
// mem_wrbits: メモリの書き込みビットマスク
// ir_ld:      IRレジスタの書き込み制御
// rs1_addr:   RS1アドレス
// rs2_addr:   RS2アドレス
// rd_addr:    RDアドレス
// rd_sel:     RDの入力選択
// rd_ld:      RDの書き込み制御
// a_ld:       Aレジスタの書き込み制御
// b_ld:       Bレジスタの書き込み制御
// a_sel:      ALUの入力1の入力選択
// b_sel:      ALUの入力2の入力選択
// imm:        即値
// alu_ctl:    ALUの機能コード
// c_ld:       Cレジスタの書き込み制御
module controller(input [3:0]	cstate,
        input [31:0]			ir,
        input [31:0] 			addr,
        input [31:0]  			alu_out,
        output    				pc_sel,
        output    				pc_ld,
        output    				mem_sel,
        output    				mem_read,
        output    				mem_write,
        output [3:0]    		mem_wrbits,
        output    				ir_ld,
        output [4:0]    		rs1_addr,
        output [4:0]    		rs2_addr,
        output [4:0]    		rd_addr,
        output [1:0]    		rd_sel,
        output    				rd_ld,
        output    				a_ld,
        output    				b_ld,
        output    				a_sel,
        output    				b_sel,
        output [31:0] 			imm,
        output [3:0]    		alu_ctl,
        output    				c_ld);

endmodule // controller
